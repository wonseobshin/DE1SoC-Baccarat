module card7seg(input [3:0] card, output[6:0] seg7);

   // your code goes here

endmodule

