module card7seg(input [3:0] SW, output [6:0] HEX0);
		
   // your code goes here
	
endmodule

